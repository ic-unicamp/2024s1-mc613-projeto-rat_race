`define VELOCIDADE_BARRA_V 40
`define VELOCIDADE_BARRA_V 40
`define ALTURA_BARRA 60
`define LARGURA_BARRA 20

  `define LIMITE_TELA_DIR 630
  `define LIMITE_TELA_ESQ 10
  `define LIMITE_TELA_CIMA 10
  `define LIMITE_TELA_BAIXO 470
  
  `define LIMITE_GOL_CIMA 180
  `define LIMITE_GOL_BAIXO 300
  
  
  
  //largura bordinhas 10
  
  //começa em 180 e termina 300 (o gol)