`define BARRA_PARADA 2'b00
`define BARRA_CIMA 2'b01
`define PORRADAO_NULL 2'b00
`define PORRADAO_INDO 2'b01
`define PORRADAO_VOLTANDO 2'b10
`define BARRA_BAIXO 2'b10
`define VELOCIDADE_BARRA_V 40
`define VELOCIDADE_PORRADAO 20
`define VELOCIDADE_BARRA_V 40
`define ALTURA_BARRA 60
`define LARGURA_BARRA 20

  `define LIMITE_TELA_DIR 640
  `define LIMITE_TELA_ESQ 0
  `define LIMITE_TELA_CIMA 0
  `define LIMITE_TELA_BAIXO 480