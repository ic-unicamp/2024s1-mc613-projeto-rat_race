module barra(
    

)


endmodule